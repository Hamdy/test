module main

fn main(){
	println("Hey")
} 